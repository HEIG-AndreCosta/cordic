--------------------------------------------------------------------------------
-- HEIG-VD
-- Haute Ecole d'Ingenerie et de Gestion du Canton de Vaud
-- School of Business and Engineering in Canton de Vaud
--------------------------------------------------------------------------------
-- REDS Institute
-- Reconfigurable Embedded Digital Systems
--------------------------------------------------------------------------------
--
-- File     : cordic_arch_pipeline.vhd
-- Author   : Yann Thoma
-- Date     : 10.04.2025
--
-- Context  : SCF lab 08
--
--------------------------------------------------------------------------------
-- Description :  Pipelined CORDIC architecture
--------------------------------------------------------------------------------
-- Dependencies : - 
--
--------------------------------------------------------------------------------
-- Modifications :
-- Ver    Date        Engineer    Comments
-- 0.1    See header  PPC         Initial version
--------------------------------------------------------------------------------

architecture pipeline of cordic is

    component cordic_pre_treatment is
        port (
                 re_i                    : in  std_logic_vector(DATASIZE - 1 downto 0);
                 im_i                    : in  std_logic_vector(DATASIZE - 1 downto 0);
                 re_o                    : out  std_logic_vector(DATASIZE - 1 downto 0);
                 im_o                    : out  std_logic_vector(DATASIZE - 1 downto 0);
                 original_quadrant_id_o  : out std_logic_vector(1 downto 0);
                 signals_exchanged_o     : out std_logic
             );
    end component;

    component cordic_iteration is
        port (
                 re_i  : in  std_logic_vector(DATASIZE - 1 downto 0);   
                 im_i  : in  std_logic_vector(DATASIZE - 1 downto 0);    
                 phi_i : in  std_logic_vector(PHI_OUTPUTSIZE - 1 downto 0);
                 re_o  : out std_logic_vector(DATASIZE - 1 downto 0);    
                 im_o  : out std_logic_vector(DATASIZE - 1 downto 0);     
                 phi_o : out std_logic_vector(PHI_OUTPUTSIZE - 1 downto 0);
                 iter_i : in std_logic_vector(3 downto 0)
             );
    end component;

    component cordic_post_treatment is
        port (
                 re_i                    : in  std_logic_vector(DATASIZE - 1 downto 0);
                 im_i                    : in  std_logic_vector(DATASIZE - 1 downto 0);
                 original_quadrant_id_i  : in std_logic_vector(1 downto 0);
                 signals_exchanged_i     : in std_logic;
                 phi_i                   : in std_logic_vector(PHI_OUTPUTSIZE - 1 downto 0);
                 amp_o       : out std_logic_vector(AMP_OUTPUTSIZE - 1 downto 0);
                 phi_o       : out std_logic_vector(PHI_OUTPUTSIZE - 1 downto 0)
             );
    end component;

    type iter_values_array_t is array (0 to 11) of std_logic_vector(DATASIZE - 1 downto 0);
    type iter_phi_array_t is array (0 to 11) of std_logic_vector(PHI_OUTPUTSIZE - 1 downto 0);
    type iter_data_valid_array_t is array (0 to 11) of std_logic;

    signal re_i_s                   : iter_values_array_t; 
    signal im_i_s                   : iter_values_array_t; 
    signal phi_i_s                  : iter_phi_array_t; 
    signal re_o_s                   : iter_values_array_t; 
    signal im_o_s                   : iter_values_array_t; 
    signal phi_o_s                  : iter_phi_array_t; 

    signal data_valid_s             : iter_data_valid_array_t;
    signal stop_s                   : iter_data_valid_array_t;
    signal original_quadrant_id_s   : std_logic_vector(1 downto 0);
    signal signals_exchanged_s      : std_logic;

    signal amp_s       :  std_logic_vector(amp_o'range);
    signal phi_s       :  std_logic_vector(phi_o'range);
    signal ready_s : std_logic;

begin
    pre_treatment: entity work.cordic_pre_treatment
    port map(
       clk_i => clk_i,
       rst_i => rst_i,
       re_i => re_i_s(0),
       im_i => im_i_s(0),
       re_o => re_o_s(0),
       im_o => re_o_s(0),
       original_quadrant_id_o => original_quadrant_id_s,
       signals_exchanged_o => signals_exchanged_s
    );

    process(clk_i)
    begin
        if rising_edge(clk_i) then
            if stop_s = '0' then
                re_i_s(1) <= re_o_s(0);
                im_i_s(1) <= re_o_s(0);
                phi_i_s(0) <= (others => '0');
                data_valid_s(0) <= ready_s and valid_i;
            end if;
        end if;
    end process;
    
    cordic_iterations: for i in 1 to 10 generate
        iteration: cordic_iteration port map (
            re_i  => re_i_s(i),   
            im_i  => im_i_s(i), 
            phi_i => phi_i_s(i - 1),
            re_o  => re_o_s(i + 1),    
            im_o  => im_o_s(i + 1),
            phi_o => phi_o_s(i),
            iter_i => std_logic_vector(to_unsigned(i + 1, 4))
        );
        process(clk_i)
        begin
            if rising_edge(clk_i) then
                if stop_s = '0' then
                    re_i_s(i + 1) <= re_o_s(i + 1);
                    re_i_s(i + 1) <= im_o_s(i + 1);
                    phi_i_s(i) <= phi_o_s(i - 1);
                    data_valid_s(i) <= data_valid_s(i - 1);
                end if;
            end if;
        end process;
    end generate;

    post_treatment: entity work.cordic_post_treatment
    port map(
       clk_i => clk_i,
       rst_i => rst_i,
       re_i => re_i_s(11),
       im_i => im_i_s(11),
       original_quadrant_id_i => original_quadrant_id_s,
       signals_exchanged_i => signals_exchanged_s,
       phi_i => phi_i_s(11),
       amp_o => amp_s,
       phi_o => phi_s
    );

    process(clk_i)
    begin
        if rising_edge(clk_i) then
            if ready_i = '1' then
                amp_o <= amp_s;
                phi_o <= phi_s;
            end if;
            valid_o <= data_valid_s(10);
        end if;
    end process;

    -- TODO: Generate stop signal for each pipeline stage
    stop_s <= data_valid_s(10) = '1' and ready_i = '0';
    ready_s <= not stop_s;
    ready_o <= ready_s;

end pipeline;
